* Vishay IRF840APBF Advanced SPICE Model
* 500 V, 8 A N-Channel MOSFET
* Extracted from datasheet 91065, Rev. C (2021)

.SUBCKT IRF840APBF D G S
* Main MOSFET (Level 3)
M1 D G S S IRF840APBF_MOD
+ L=1u W=1u 
+ M=1 

* Gate Resistance
RG G G1 0.7  ; Gate input resistance (typ. 0.7 Ω, max. 3.7 Ω)

* Drain-Source Resistances
RD D D1 0.0425 ; RDS(on)/2 (typ. 0.085 Ω @ VGS=10 V, ID=4.8 A)
RS S S1 0.0425

* Capacitances (from Ciss, Coss, Crss)
CGS G S 1.8n  ; Ciss - Crss = 1018 pF - 8 pF ≈ 1.8 nF
CGD G D 100p   ; Crss = 8 pF (typ.)
CDS D S 155p   ; Coss - Cgd = 155 pF - 8 pF ≈ 155 pF

* Body Diode
D1 S D IRF840APBF_DIODE

* Models
.MODEL IRF840APBF_MOD NMOS (
+ LEVEL=3 VTO=4 KP=10 LAMBDA=0.01 
+ RS=0.0425 RD=0.0425 RDS=1E6 
+ IS=1E-12 N=1.5 TT=422n 
+ CGSO=1.8n CGDO=100p CGBO=1p 
+ TOX=100n NSUB=1E15 UO=600 
+ KF=1E-28 AF=1 FC=0.5
)

.MODEL IRF840APBF_DIODE D (
+ IS=1E-11 RS=0.0425 N=1.5 TT=422n 
+ CJO=155p VJ=0.8 M=0.5
)

* Thermal Parameters (RthJC = 1.0 °C/W)
.THERMAL RTHJC=1.0 RTHCS=0.5

.ENDS IRF840APBF