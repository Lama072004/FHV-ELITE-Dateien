* Nexperia PHP79NQ08LT - Enhanced Model
.SUBCKT PHP79NQ08LT D G S
M1 D G S S NXP_NMOS L=1u W=500u
.MODEL NXP_NMOS NMOS LEVEL=1
+ VTO=1.5
+ KP=120e-6
+ LAMBDA=0.01
+ RDS=0.015
+ CGSO=0.8n CGDO=0.3n
+ CBD=300p CBS=300p
+ IS=1e-9 PB=0.8 MJ=0.5
D1 S D Dbody
.MODEL Dbody D IS=1e-9 N=1 TT=100n RS=0.02
.ENDS PHP79NQ08LT
