* Nexperia PHP79NQ08LT Advanced SPICE Model
* 75 V, 73 A Logic-Level N-Channel MOSFET
* Extracted from datasheet Rev. 03 (2010)

.SUBCKT PHP79NQ08LT D G S
* Main MOSFET (Level 3)
M1 D G S S PHP79NQ08LT_MOD
+ L=1u W=1u 
+ M=1 

* Gate Resistance
RG G G1 1.0  ; Estimated (datasheet lacks Rg)

* Drain-Source Resistances
RD D D1 0.007 ; RDS(on)/2 (typ. 14 mΩ @ VGS=10 V, ID=25 A)
RS S S1 0.007

* Capacitances (from Ciss, Coss, Crss)
CGS G S 2.9n  ; Ciss - Crss = 3026 pF - 140 pF ≈ 2.9 nF
CGD G D 140p   ; Crss = 140 pF (typ.)
CDS D S 161p   ; Coss - Cgd = 301 pF - 140 pF ≈ 161 pF

* Body Diode
D1 S D PHP79NQ08LT_DIODE

* Models
.MODEL PHP79NQ08LT_MOD NMOS (
+ LEVEL=3 VTO=1.5 KP=30 LAMBDA=0.02 
+ RS=0.007 RD=0.007 RDS=1E6 
+ IS=1E-12 N=1.5 TT=90n 
+ CGSO=2.9n CGDO=140p CGBO=1p 
+ TOX=100n NSUB=1E15 UO=700 
+ KF=1E-28 AF=1 FC=0.5
)

.MODEL PHP79NQ08LT_DIODE D (
+ IS=1E-11 RS=0.007 N=1.5 TT=90n 
+ CJO=161p VJ=0.8 M=0.5
)

* Thermal Parameters (RthJC = 0.95 K/W)
.THERMAL RTHJC=0.95 RTHCS=0.5

.ENDS PHP79NQ08LT