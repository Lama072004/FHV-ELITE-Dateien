* Vishay IRF840A - Enhanced Model
.SUBCKT IRF840A D G S
M1 D G S S VISHAY_NMOS L=1u W=300u
.MODEL VISHAY_NMOS NMOS LEVEL=1
+ VTO=3.0
+ KP=45e-6
+ LAMBDA=0.01
+ RDS=0.85
+ CGSO=1.2n CGDO=0.6n
+ CBD=150p CBS=150p
+ IS=1e-9 PB=0.8 MJ=0.5
D1 S D Dbody
.MODEL Dbody D IS=1e-9 N=1 TT=422n RS=0.02
.ENDS IRF840A
